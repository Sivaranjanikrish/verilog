module constantio(in,out);
	output out;
	input in;
	assign out=in;
endmodule
