module BCDto7segdf(bcd,seg);
	output[6:0]seg;
	input[3:0]bcd;
  assign seg=
	  (bcd == 4'b0000) ? 7'b1111110 :  
          (bcd == 4'b0001) ? 7'b0110000 :  
          (bcd == 4'b0010) ? 7'b1101101 :  
	  (bcd == 4'b0011) ? 7'b1111001 :  
          (bcd == 4'b0100) ? 7'b0110011 :  
          (bcd == 4'b0101) ? 7'b1011011 :  
         (bcd == 4'b0110) ? 7'b1011111 :  
         (bcd == 4'b0111) ? 7'b1110000 :
    (bcd == 4'b1000) ? 7'b1111111 :  
       (bcd == 4'b1001) ? 7'b1111011 :
	7'b0000000;
endmodule
