module constant1(output out);
	assign out=1'b1;
endmodule
