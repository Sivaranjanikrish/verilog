module constant_0(output out);
	assign out=1'b0;
endmodule
